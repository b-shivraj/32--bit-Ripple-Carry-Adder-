module RCA_32 (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire c1;
 wire c2;
 wire c3;
 wire \M0/c1 ;
 wire \M0/M0/c1 ;
 wire \M0/M0/c2 ;
 wire \M0/M0/c3 ;
 wire \M0/M0/M0/_0_ ;
 wire \M0/M0/M0/_1_ ;
 wire \M0/M0/M0/_2_ ;
 wire \M0/M0/M0/_3_ ;
 wire \M0/M0/M1/_0_ ;
 wire \M0/M0/M1/_1_ ;
 wire \M0/M0/M1/_2_ ;
 wire \M0/M0/M1/_3_ ;
 wire \M0/M0/M2/_0_ ;
 wire \M0/M0/M2/_1_ ;
 wire \M0/M0/M2/_2_ ;
 wire \M0/M0/M2/_3_ ;
 wire \M0/M0/M3/_0_ ;
 wire \M0/M0/M3/_1_ ;
 wire \M0/M0/M3/_2_ ;
 wire \M0/M0/M3/_3_ ;
 wire \M0/M1/c1 ;
 wire \M0/M1/c2 ;
 wire \M0/M1/c3 ;
 wire \M0/M1/M0/_0_ ;
 wire \M0/M1/M0/_1_ ;
 wire \M0/M1/M0/_2_ ;
 wire \M0/M1/M0/_3_ ;
 wire \M0/M1/M1/_0_ ;
 wire \M0/M1/M1/_1_ ;
 wire \M0/M1/M1/_2_ ;
 wire \M0/M1/M1/_3_ ;
 wire \M0/M1/M2/_0_ ;
 wire \M0/M1/M2/_1_ ;
 wire \M0/M1/M2/_2_ ;
 wire \M0/M1/M2/_3_ ;
 wire \M0/M1/M3/_0_ ;
 wire \M0/M1/M3/_1_ ;
 wire \M0/M1/M3/_2_ ;
 wire \M0/M1/M3/_3_ ;
 wire \M1/c1 ;
 wire \M1/M0/c1 ;
 wire \M1/M0/c2 ;
 wire \M1/M0/c3 ;
 wire \M1/M0/M0/_0_ ;
 wire \M1/M0/M0/_1_ ;
 wire \M1/M0/M0/_2_ ;
 wire \M1/M0/M0/_3_ ;
 wire \M1/M0/M1/_0_ ;
 wire \M1/M0/M1/_1_ ;
 wire \M1/M0/M1/_2_ ;
 wire \M1/M0/M1/_3_ ;
 wire \M1/M0/M2/_0_ ;
 wire \M1/M0/M2/_1_ ;
 wire \M1/M0/M2/_2_ ;
 wire \M1/M0/M2/_3_ ;
 wire \M1/M0/M3/_0_ ;
 wire \M1/M0/M3/_1_ ;
 wire \M1/M0/M3/_2_ ;
 wire \M1/M0/M3/_3_ ;
 wire \M1/M1/c1 ;
 wire \M1/M1/c2 ;
 wire \M1/M1/c3 ;
 wire \M1/M1/M0/_0_ ;
 wire \M1/M1/M0/_1_ ;
 wire \M1/M1/M0/_2_ ;
 wire \M1/M1/M0/_3_ ;
 wire \M1/M1/M1/_0_ ;
 wire \M1/M1/M1/_1_ ;
 wire \M1/M1/M1/_2_ ;
 wire \M1/M1/M1/_3_ ;
 wire \M1/M1/M2/_0_ ;
 wire \M1/M1/M2/_1_ ;
 wire \M1/M1/M2/_2_ ;
 wire \M1/M1/M2/_3_ ;
 wire \M1/M1/M3/_0_ ;
 wire \M1/M1/M3/_1_ ;
 wire \M1/M1/M3/_2_ ;
 wire \M1/M1/M3/_3_ ;
 wire \M2/c1 ;
 wire \M2/M0/c1 ;
 wire \M2/M0/c2 ;
 wire \M2/M0/c3 ;
 wire \M2/M0/M0/_0_ ;
 wire \M2/M0/M0/_1_ ;
 wire \M2/M0/M0/_2_ ;
 wire \M2/M0/M0/_3_ ;
 wire \M2/M0/M1/_0_ ;
 wire \M2/M0/M1/_1_ ;
 wire \M2/M0/M1/_2_ ;
 wire \M2/M0/M1/_3_ ;
 wire \M2/M0/M2/_0_ ;
 wire \M2/M0/M2/_1_ ;
 wire \M2/M0/M2/_2_ ;
 wire \M2/M0/M2/_3_ ;
 wire \M2/M0/M3/_0_ ;
 wire \M2/M0/M3/_1_ ;
 wire \M2/M0/M3/_2_ ;
 wire \M2/M0/M3/_3_ ;
 wire \M2/M1/c1 ;
 wire \M2/M1/c2 ;
 wire \M2/M1/c3 ;
 wire \M2/M1/M0/_0_ ;
 wire \M2/M1/M0/_1_ ;
 wire \M2/M1/M0/_2_ ;
 wire \M2/M1/M0/_3_ ;
 wire \M2/M1/M1/_0_ ;
 wire \M2/M1/M1/_1_ ;
 wire \M2/M1/M1/_2_ ;
 wire \M2/M1/M1/_3_ ;
 wire \M2/M1/M2/_0_ ;
 wire \M2/M1/M2/_1_ ;
 wire \M2/M1/M2/_2_ ;
 wire \M2/M1/M2/_3_ ;
 wire \M2/M1/M3/_0_ ;
 wire \M2/M1/M3/_1_ ;
 wire \M2/M1/M3/_2_ ;
 wire \M2/M1/M3/_3_ ;
 wire \M3/c1 ;
 wire \M3/M0/c1 ;
 wire \M3/M0/c2 ;
 wire \M3/M0/c3 ;
 wire \M3/M0/M0/_0_ ;
 wire \M3/M0/M0/_1_ ;
 wire \M3/M0/M0/_2_ ;
 wire \M3/M0/M0/_3_ ;
 wire \M3/M0/M1/_0_ ;
 wire \M3/M0/M1/_1_ ;
 wire \M3/M0/M1/_2_ ;
 wire \M3/M0/M1/_3_ ;
 wire \M3/M0/M2/_0_ ;
 wire \M3/M0/M2/_1_ ;
 wire \M3/M0/M2/_2_ ;
 wire \M3/M0/M2/_3_ ;
 wire \M3/M0/M3/_0_ ;
 wire \M3/M0/M3/_1_ ;
 wire \M3/M0/M3/_2_ ;
 wire \M3/M0/M3/_3_ ;
 wire \M3/M1/c1 ;
 wire \M3/M1/c2 ;
 wire \M3/M1/c3 ;
 wire \M3/M1/M0/_0_ ;
 wire \M3/M1/M0/_1_ ;
 wire \M3/M1/M0/_2_ ;
 wire \M3/M1/M0/_3_ ;
 wire \M3/M1/M1/_0_ ;
 wire \M3/M1/M1/_1_ ;
 wire \M3/M1/M1/_2_ ;
 wire \M3/M1/M1/_3_ ;
 wire \M3/M1/M2/_0_ ;
 wire \M3/M1/M2/_1_ ;
 wire \M3/M1/M2/_2_ ;
 wire \M3/M1/M2/_3_ ;
 wire \M3/M1/M3/_0_ ;
 wire \M3/M1/M3/_1_ ;
 wire \M3/M1/M3/_2_ ;
 wire \M3/M1/M3/_3_ ;

 INV_X1 \M0/M0/M0/_4_  (.A(cin),
    .ZN(\M0/M0/M0/_0_ ));
 NAND2_X1 \M0/M0/M0/_5_  (.A1(a[0]),
    .A2(b[0]),
    .ZN(\M0/M0/M0/_1_ ));
 NOR2_X1 \M0/M0/M0/_6_  (.A1(a[0]),
    .A2(b[0]),
    .ZN(\M0/M0/M0/_2_ ));
 XOR2_X1 \M0/M0/M0/_7_  (.A(a[0]),
    .B(b[0]),
    .Z(\M0/M0/M0/_3_ ));
 OAI21_X1 \M0/M0/M0/_8_  (.A(\M0/M0/M0/_1_ ),
    .B1(\M0/M0/M0/_2_ ),
    .B2(\M0/M0/M0/_0_ ),
    .ZN(\M0/M0/c1 ));
 XNOR2_X1 \M0/M0/M0/_9_  (.A(\M0/M0/M0/_0_ ),
    .B(\M0/M0/M0/_3_ ),
    .ZN(sum[0]));
 INV_X1 \M0/M0/M1/_4_  (.A(\M0/M0/c1 ),
    .ZN(\M0/M0/M1/_0_ ));
 NAND2_X1 \M0/M0/M1/_5_  (.A1(a[1]),
    .A2(b[1]),
    .ZN(\M0/M0/M1/_1_ ));
 NOR2_X1 \M0/M0/M1/_6_  (.A1(a[1]),
    .A2(b[1]),
    .ZN(\M0/M0/M1/_2_ ));
 XOR2_X1 \M0/M0/M1/_7_  (.A(a[1]),
    .B(b[1]),
    .Z(\M0/M0/M1/_3_ ));
 OAI21_X1 \M0/M0/M1/_8_  (.A(\M0/M0/M1/_1_ ),
    .B1(\M0/M0/M1/_2_ ),
    .B2(\M0/M0/M1/_0_ ),
    .ZN(\M0/M0/c2 ));
 XNOR2_X1 \M0/M0/M1/_9_  (.A(\M0/M0/M1/_0_ ),
    .B(\M0/M0/M1/_3_ ),
    .ZN(sum[1]));
 INV_X1 \M0/M0/M2/_4_  (.A(\M0/M0/c2 ),
    .ZN(\M0/M0/M2/_0_ ));
 NAND2_X1 \M0/M0/M2/_5_  (.A1(a[2]),
    .A2(b[2]),
    .ZN(\M0/M0/M2/_1_ ));
 NOR2_X1 \M0/M0/M2/_6_  (.A1(a[2]),
    .A2(b[2]),
    .ZN(\M0/M0/M2/_2_ ));
 XOR2_X1 \M0/M0/M2/_7_  (.A(a[2]),
    .B(b[2]),
    .Z(\M0/M0/M2/_3_ ));
 OAI21_X1 \M0/M0/M2/_8_  (.A(\M0/M0/M2/_1_ ),
    .B1(\M0/M0/M2/_2_ ),
    .B2(\M0/M0/M2/_0_ ),
    .ZN(\M0/M0/c3 ));
 XNOR2_X1 \M0/M0/M2/_9_  (.A(\M0/M0/M2/_0_ ),
    .B(\M0/M0/M2/_3_ ),
    .ZN(sum[2]));
 INV_X1 \M0/M0/M3/_4_  (.A(\M0/M0/c3 ),
    .ZN(\M0/M0/M3/_0_ ));
 NAND2_X1 \M0/M0/M3/_5_  (.A1(a[3]),
    .A2(b[3]),
    .ZN(\M0/M0/M3/_1_ ));
 NOR2_X1 \M0/M0/M3/_6_  (.A1(a[3]),
    .A2(b[3]),
    .ZN(\M0/M0/M3/_2_ ));
 XOR2_X1 \M0/M0/M3/_7_  (.A(a[3]),
    .B(b[3]),
    .Z(\M0/M0/M3/_3_ ));
 OAI21_X1 \M0/M0/M3/_8_  (.A(\M0/M0/M3/_1_ ),
    .B1(\M0/M0/M3/_2_ ),
    .B2(\M0/M0/M3/_0_ ),
    .ZN(\M0/c1 ));
 XNOR2_X1 \M0/M0/M3/_9_  (.A(\M0/M0/M3/_0_ ),
    .B(\M0/M0/M3/_3_ ),
    .ZN(sum[3]));
 INV_X1 \M0/M1/M0/_4_  (.A(\M0/c1 ),
    .ZN(\M0/M1/M0/_0_ ));
 NAND2_X1 \M0/M1/M0/_5_  (.A1(a[4]),
    .A2(b[4]),
    .ZN(\M0/M1/M0/_1_ ));
 NOR2_X1 \M0/M1/M0/_6_  (.A1(a[4]),
    .A2(b[4]),
    .ZN(\M0/M1/M0/_2_ ));
 XOR2_X1 \M0/M1/M0/_7_  (.A(a[4]),
    .B(b[4]),
    .Z(\M0/M1/M0/_3_ ));
 OAI21_X1 \M0/M1/M0/_8_  (.A(\M0/M1/M0/_1_ ),
    .B1(\M0/M1/M0/_2_ ),
    .B2(\M0/M1/M0/_0_ ),
    .ZN(\M0/M1/c1 ));
 XNOR2_X1 \M0/M1/M0/_9_  (.A(\M0/M1/M0/_0_ ),
    .B(\M0/M1/M0/_3_ ),
    .ZN(sum[4]));
 INV_X1 \M0/M1/M1/_4_  (.A(\M0/M1/c1 ),
    .ZN(\M0/M1/M1/_0_ ));
 NAND2_X1 \M0/M1/M1/_5_  (.A1(a[5]),
    .A2(b[5]),
    .ZN(\M0/M1/M1/_1_ ));
 NOR2_X1 \M0/M1/M1/_6_  (.A1(a[5]),
    .A2(b[5]),
    .ZN(\M0/M1/M1/_2_ ));
 XOR2_X1 \M0/M1/M1/_7_  (.A(a[5]),
    .B(b[5]),
    .Z(\M0/M1/M1/_3_ ));
 OAI21_X1 \M0/M1/M1/_8_  (.A(\M0/M1/M1/_1_ ),
    .B1(\M0/M1/M1/_2_ ),
    .B2(\M0/M1/M1/_0_ ),
    .ZN(\M0/M1/c2 ));
 XNOR2_X1 \M0/M1/M1/_9_  (.A(\M0/M1/M1/_0_ ),
    .B(\M0/M1/M1/_3_ ),
    .ZN(sum[5]));
 INV_X1 \M0/M1/M2/_4_  (.A(\M0/M1/c2 ),
    .ZN(\M0/M1/M2/_0_ ));
 NAND2_X1 \M0/M1/M2/_5_  (.A1(a[6]),
    .A2(b[6]),
    .ZN(\M0/M1/M2/_1_ ));
 NOR2_X1 \M0/M1/M2/_6_  (.A1(a[6]),
    .A2(b[6]),
    .ZN(\M0/M1/M2/_2_ ));
 XOR2_X1 \M0/M1/M2/_7_  (.A(a[6]),
    .B(b[6]),
    .Z(\M0/M1/M2/_3_ ));
 OAI21_X1 \M0/M1/M2/_8_  (.A(\M0/M1/M2/_1_ ),
    .B1(\M0/M1/M2/_2_ ),
    .B2(\M0/M1/M2/_0_ ),
    .ZN(\M0/M1/c3 ));
 XNOR2_X1 \M0/M1/M2/_9_  (.A(\M0/M1/M2/_0_ ),
    .B(\M0/M1/M2/_3_ ),
    .ZN(sum[6]));
 INV_X1 \M0/M1/M3/_4_  (.A(\M0/M1/c3 ),
    .ZN(\M0/M1/M3/_0_ ));
 NAND2_X1 \M0/M1/M3/_5_  (.A1(a[7]),
    .A2(b[7]),
    .ZN(\M0/M1/M3/_1_ ));
 NOR2_X1 \M0/M1/M3/_6_  (.A1(a[7]),
    .A2(b[7]),
    .ZN(\M0/M1/M3/_2_ ));
 XOR2_X1 \M0/M1/M3/_7_  (.A(a[7]),
    .B(b[7]),
    .Z(\M0/M1/M3/_3_ ));
 OAI21_X1 \M0/M1/M3/_8_  (.A(\M0/M1/M3/_1_ ),
    .B1(\M0/M1/M3/_2_ ),
    .B2(\M0/M1/M3/_0_ ),
    .ZN(c1));
 XNOR2_X1 \M0/M1/M3/_9_  (.A(\M0/M1/M3/_0_ ),
    .B(\M0/M1/M3/_3_ ),
    .ZN(sum[7]));
 INV_X1 \M1/M0/M0/_4_  (.A(c1),
    .ZN(\M1/M0/M0/_0_ ));
 NAND2_X1 \M1/M0/M0/_5_  (.A1(a[8]),
    .A2(b[8]),
    .ZN(\M1/M0/M0/_1_ ));
 NOR2_X1 \M1/M0/M0/_6_  (.A1(a[8]),
    .A2(b[8]),
    .ZN(\M1/M0/M0/_2_ ));
 XOR2_X1 \M1/M0/M0/_7_  (.A(a[8]),
    .B(b[8]),
    .Z(\M1/M0/M0/_3_ ));
 OAI21_X1 \M1/M0/M0/_8_  (.A(\M1/M0/M0/_1_ ),
    .B1(\M1/M0/M0/_2_ ),
    .B2(\M1/M0/M0/_0_ ),
    .ZN(\M1/M0/c1 ));
 XNOR2_X1 \M1/M0/M0/_9_  (.A(\M1/M0/M0/_0_ ),
    .B(\M1/M0/M0/_3_ ),
    .ZN(sum[8]));
 INV_X1 \M1/M0/M1/_4_  (.A(\M1/M0/c1 ),
    .ZN(\M1/M0/M1/_0_ ));
 NAND2_X1 \M1/M0/M1/_5_  (.A1(a[9]),
    .A2(b[9]),
    .ZN(\M1/M0/M1/_1_ ));
 NOR2_X1 \M1/M0/M1/_6_  (.A1(a[9]),
    .A2(b[9]),
    .ZN(\M1/M0/M1/_2_ ));
 XOR2_X1 \M1/M0/M1/_7_  (.A(a[9]),
    .B(b[9]),
    .Z(\M1/M0/M1/_3_ ));
 OAI21_X1 \M1/M0/M1/_8_  (.A(\M1/M0/M1/_1_ ),
    .B1(\M1/M0/M1/_2_ ),
    .B2(\M1/M0/M1/_0_ ),
    .ZN(\M1/M0/c2 ));
 XNOR2_X1 \M1/M0/M1/_9_  (.A(\M1/M0/M1/_0_ ),
    .B(\M1/M0/M1/_3_ ),
    .ZN(sum[9]));
 INV_X1 \M1/M0/M2/_4_  (.A(\M1/M0/c2 ),
    .ZN(\M1/M0/M2/_0_ ));
 NAND2_X1 \M1/M0/M2/_5_  (.A1(a[10]),
    .A2(b[10]),
    .ZN(\M1/M0/M2/_1_ ));
 NOR2_X1 \M1/M0/M2/_6_  (.A1(a[10]),
    .A2(b[10]),
    .ZN(\M1/M0/M2/_2_ ));
 XOR2_X1 \M1/M0/M2/_7_  (.A(a[10]),
    .B(b[10]),
    .Z(\M1/M0/M2/_3_ ));
 OAI21_X1 \M1/M0/M2/_8_  (.A(\M1/M0/M2/_1_ ),
    .B1(\M1/M0/M2/_2_ ),
    .B2(\M1/M0/M2/_0_ ),
    .ZN(\M1/M0/c3 ));
 XNOR2_X1 \M1/M0/M2/_9_  (.A(\M1/M0/M2/_0_ ),
    .B(\M1/M0/M2/_3_ ),
    .ZN(sum[10]));
 INV_X1 \M1/M0/M3/_4_  (.A(\M1/M0/c3 ),
    .ZN(\M1/M0/M3/_0_ ));
 NAND2_X1 \M1/M0/M3/_5_  (.A1(a[11]),
    .A2(b[11]),
    .ZN(\M1/M0/M3/_1_ ));
 NOR2_X1 \M1/M0/M3/_6_  (.A1(a[11]),
    .A2(b[11]),
    .ZN(\M1/M0/M3/_2_ ));
 XOR2_X1 \M1/M0/M3/_7_  (.A(a[11]),
    .B(b[11]),
    .Z(\M1/M0/M3/_3_ ));
 OAI21_X1 \M1/M0/M3/_8_  (.A(\M1/M0/M3/_1_ ),
    .B1(\M1/M0/M3/_2_ ),
    .B2(\M1/M0/M3/_0_ ),
    .ZN(\M1/c1 ));
 XNOR2_X1 \M1/M0/M3/_9_  (.A(\M1/M0/M3/_0_ ),
    .B(\M1/M0/M3/_3_ ),
    .ZN(sum[11]));
 INV_X1 \M1/M1/M0/_4_  (.A(\M1/c1 ),
    .ZN(\M1/M1/M0/_0_ ));
 NAND2_X1 \M1/M1/M0/_5_  (.A1(a[12]),
    .A2(b[12]),
    .ZN(\M1/M1/M0/_1_ ));
 NOR2_X1 \M1/M1/M0/_6_  (.A1(a[12]),
    .A2(b[12]),
    .ZN(\M1/M1/M0/_2_ ));
 XOR2_X1 \M1/M1/M0/_7_  (.A(a[12]),
    .B(b[12]),
    .Z(\M1/M1/M0/_3_ ));
 OAI21_X1 \M1/M1/M0/_8_  (.A(\M1/M1/M0/_1_ ),
    .B1(\M1/M1/M0/_2_ ),
    .B2(\M1/M1/M0/_0_ ),
    .ZN(\M1/M1/c1 ));
 XNOR2_X1 \M1/M1/M0/_9_  (.A(\M1/M1/M0/_0_ ),
    .B(\M1/M1/M0/_3_ ),
    .ZN(sum[12]));
 INV_X1 \M1/M1/M1/_4_  (.A(\M1/M1/c1 ),
    .ZN(\M1/M1/M1/_0_ ));
 NAND2_X1 \M1/M1/M1/_5_  (.A1(a[13]),
    .A2(b[13]),
    .ZN(\M1/M1/M1/_1_ ));
 NOR2_X1 \M1/M1/M1/_6_  (.A1(a[13]),
    .A2(b[13]),
    .ZN(\M1/M1/M1/_2_ ));
 XOR2_X1 \M1/M1/M1/_7_  (.A(a[13]),
    .B(b[13]),
    .Z(\M1/M1/M1/_3_ ));
 OAI21_X1 \M1/M1/M1/_8_  (.A(\M1/M1/M1/_1_ ),
    .B1(\M1/M1/M1/_2_ ),
    .B2(\M1/M1/M1/_0_ ),
    .ZN(\M1/M1/c2 ));
 XNOR2_X1 \M1/M1/M1/_9_  (.A(\M1/M1/M1/_0_ ),
    .B(\M1/M1/M1/_3_ ),
    .ZN(sum[13]));
 INV_X1 \M1/M1/M2/_4_  (.A(\M1/M1/c2 ),
    .ZN(\M1/M1/M2/_0_ ));
 NAND2_X1 \M1/M1/M2/_5_  (.A1(a[14]),
    .A2(b[14]),
    .ZN(\M1/M1/M2/_1_ ));
 NOR2_X1 \M1/M1/M2/_6_  (.A1(a[14]),
    .A2(b[14]),
    .ZN(\M1/M1/M2/_2_ ));
 XOR2_X1 \M1/M1/M2/_7_  (.A(a[14]),
    .B(b[14]),
    .Z(\M1/M1/M2/_3_ ));
 OAI21_X1 \M1/M1/M2/_8_  (.A(\M1/M1/M2/_1_ ),
    .B1(\M1/M1/M2/_2_ ),
    .B2(\M1/M1/M2/_0_ ),
    .ZN(\M1/M1/c3 ));
 XNOR2_X1 \M1/M1/M2/_9_  (.A(\M1/M1/M2/_0_ ),
    .B(\M1/M1/M2/_3_ ),
    .ZN(sum[14]));
 INV_X1 \M1/M1/M3/_4_  (.A(\M1/M1/c3 ),
    .ZN(\M1/M1/M3/_0_ ));
 NAND2_X1 \M1/M1/M3/_5_  (.A1(a[15]),
    .A2(b[15]),
    .ZN(\M1/M1/M3/_1_ ));
 NOR2_X1 \M1/M1/M3/_6_  (.A1(a[15]),
    .A2(b[15]),
    .ZN(\M1/M1/M3/_2_ ));
 XOR2_X1 \M1/M1/M3/_7_  (.A(a[15]),
    .B(b[15]),
    .Z(\M1/M1/M3/_3_ ));
 OAI21_X1 \M1/M1/M3/_8_  (.A(\M1/M1/M3/_1_ ),
    .B1(\M1/M1/M3/_2_ ),
    .B2(\M1/M1/M3/_0_ ),
    .ZN(c2));
 XNOR2_X1 \M1/M1/M3/_9_  (.A(\M1/M1/M3/_0_ ),
    .B(\M1/M1/M3/_3_ ),
    .ZN(sum[15]));
 INV_X1 \M2/M0/M0/_4_  (.A(c2),
    .ZN(\M2/M0/M0/_0_ ));
 NAND2_X1 \M2/M0/M0/_5_  (.A1(a[16]),
    .A2(b[16]),
    .ZN(\M2/M0/M0/_1_ ));
 NOR2_X1 \M2/M0/M0/_6_  (.A1(a[16]),
    .A2(b[16]),
    .ZN(\M2/M0/M0/_2_ ));
 XOR2_X1 \M2/M0/M0/_7_  (.A(a[16]),
    .B(b[16]),
    .Z(\M2/M0/M0/_3_ ));
 OAI21_X1 \M2/M0/M0/_8_  (.A(\M2/M0/M0/_1_ ),
    .B1(\M2/M0/M0/_2_ ),
    .B2(\M2/M0/M0/_0_ ),
    .ZN(\M2/M0/c1 ));
 XNOR2_X1 \M2/M0/M0/_9_  (.A(\M2/M0/M0/_0_ ),
    .B(\M2/M0/M0/_3_ ),
    .ZN(sum[16]));
 INV_X1 \M2/M0/M1/_4_  (.A(\M2/M0/c1 ),
    .ZN(\M2/M0/M1/_0_ ));
 NAND2_X1 \M2/M0/M1/_5_  (.A1(a[17]),
    .A2(b[17]),
    .ZN(\M2/M0/M1/_1_ ));
 NOR2_X1 \M2/M0/M1/_6_  (.A1(a[17]),
    .A2(b[17]),
    .ZN(\M2/M0/M1/_2_ ));
 XOR2_X1 \M2/M0/M1/_7_  (.A(a[17]),
    .B(b[17]),
    .Z(\M2/M0/M1/_3_ ));
 OAI21_X1 \M2/M0/M1/_8_  (.A(\M2/M0/M1/_1_ ),
    .B1(\M2/M0/M1/_2_ ),
    .B2(\M2/M0/M1/_0_ ),
    .ZN(\M2/M0/c2 ));
 XNOR2_X1 \M2/M0/M1/_9_  (.A(\M2/M0/M1/_0_ ),
    .B(\M2/M0/M1/_3_ ),
    .ZN(sum[17]));
 INV_X1 \M2/M0/M2/_4_  (.A(\M2/M0/c2 ),
    .ZN(\M2/M0/M2/_0_ ));
 NAND2_X1 \M2/M0/M2/_5_  (.A1(a[18]),
    .A2(b[18]),
    .ZN(\M2/M0/M2/_1_ ));
 NOR2_X1 \M2/M0/M2/_6_  (.A1(a[18]),
    .A2(b[18]),
    .ZN(\M2/M0/M2/_2_ ));
 XOR2_X1 \M2/M0/M2/_7_  (.A(a[18]),
    .B(b[18]),
    .Z(\M2/M0/M2/_3_ ));
 OAI21_X1 \M2/M0/M2/_8_  (.A(\M2/M0/M2/_1_ ),
    .B1(\M2/M0/M2/_2_ ),
    .B2(\M2/M0/M2/_0_ ),
    .ZN(\M2/M0/c3 ));
 XNOR2_X1 \M2/M0/M2/_9_  (.A(\M2/M0/M2/_0_ ),
    .B(\M2/M0/M2/_3_ ),
    .ZN(sum[18]));
 INV_X1 \M2/M0/M3/_4_  (.A(\M2/M0/c3 ),
    .ZN(\M2/M0/M3/_0_ ));
 NAND2_X1 \M2/M0/M3/_5_  (.A1(a[19]),
    .A2(b[19]),
    .ZN(\M2/M0/M3/_1_ ));
 NOR2_X1 \M2/M0/M3/_6_  (.A1(a[19]),
    .A2(b[19]),
    .ZN(\M2/M0/M3/_2_ ));
 XOR2_X1 \M2/M0/M3/_7_  (.A(a[19]),
    .B(b[19]),
    .Z(\M2/M0/M3/_3_ ));
 OAI21_X1 \M2/M0/M3/_8_  (.A(\M2/M0/M3/_1_ ),
    .B1(\M2/M0/M3/_2_ ),
    .B2(\M2/M0/M3/_0_ ),
    .ZN(\M2/c1 ));
 XNOR2_X1 \M2/M0/M3/_9_  (.A(\M2/M0/M3/_0_ ),
    .B(\M2/M0/M3/_3_ ),
    .ZN(sum[19]));
 INV_X1 \M2/M1/M0/_4_  (.A(\M2/c1 ),
    .ZN(\M2/M1/M0/_0_ ));
 NAND2_X1 \M2/M1/M0/_5_  (.A1(a[20]),
    .A2(b[20]),
    .ZN(\M2/M1/M0/_1_ ));
 NOR2_X1 \M2/M1/M0/_6_  (.A1(a[20]),
    .A2(b[20]),
    .ZN(\M2/M1/M0/_2_ ));
 XOR2_X1 \M2/M1/M0/_7_  (.A(a[20]),
    .B(b[20]),
    .Z(\M2/M1/M0/_3_ ));
 OAI21_X1 \M2/M1/M0/_8_  (.A(\M2/M1/M0/_1_ ),
    .B1(\M2/M1/M0/_2_ ),
    .B2(\M2/M1/M0/_0_ ),
    .ZN(\M2/M1/c1 ));
 XNOR2_X1 \M2/M1/M0/_9_  (.A(\M2/M1/M0/_0_ ),
    .B(\M2/M1/M0/_3_ ),
    .ZN(sum[20]));
 INV_X1 \M2/M1/M1/_4_  (.A(\M2/M1/c1 ),
    .ZN(\M2/M1/M1/_0_ ));
 NAND2_X1 \M2/M1/M1/_5_  (.A1(a[21]),
    .A2(b[21]),
    .ZN(\M2/M1/M1/_1_ ));
 NOR2_X1 \M2/M1/M1/_6_  (.A1(a[21]),
    .A2(b[21]),
    .ZN(\M2/M1/M1/_2_ ));
 XOR2_X1 \M2/M1/M1/_7_  (.A(a[21]),
    .B(b[21]),
    .Z(\M2/M1/M1/_3_ ));
 OAI21_X1 \M2/M1/M1/_8_  (.A(\M2/M1/M1/_1_ ),
    .B1(\M2/M1/M1/_2_ ),
    .B2(\M2/M1/M1/_0_ ),
    .ZN(\M2/M1/c2 ));
 XNOR2_X1 \M2/M1/M1/_9_  (.A(\M2/M1/M1/_0_ ),
    .B(\M2/M1/M1/_3_ ),
    .ZN(sum[21]));
 INV_X1 \M2/M1/M2/_4_  (.A(\M2/M1/c2 ),
    .ZN(\M2/M1/M2/_0_ ));
 NAND2_X1 \M2/M1/M2/_5_  (.A1(a[22]),
    .A2(b[22]),
    .ZN(\M2/M1/M2/_1_ ));
 NOR2_X1 \M2/M1/M2/_6_  (.A1(a[22]),
    .A2(b[22]),
    .ZN(\M2/M1/M2/_2_ ));
 XOR2_X1 \M2/M1/M2/_7_  (.A(a[22]),
    .B(b[22]),
    .Z(\M2/M1/M2/_3_ ));
 OAI21_X1 \M2/M1/M2/_8_  (.A(\M2/M1/M2/_1_ ),
    .B1(\M2/M1/M2/_2_ ),
    .B2(\M2/M1/M2/_0_ ),
    .ZN(\M2/M1/c3 ));
 XNOR2_X1 \M2/M1/M2/_9_  (.A(\M2/M1/M2/_0_ ),
    .B(\M2/M1/M2/_3_ ),
    .ZN(sum[22]));
 INV_X1 \M2/M1/M3/_4_  (.A(\M2/M1/c3 ),
    .ZN(\M2/M1/M3/_0_ ));
 NAND2_X1 \M2/M1/M3/_5_  (.A1(a[23]),
    .A2(b[23]),
    .ZN(\M2/M1/M3/_1_ ));
 NOR2_X1 \M2/M1/M3/_6_  (.A1(a[23]),
    .A2(b[23]),
    .ZN(\M2/M1/M3/_2_ ));
 XOR2_X1 \M2/M1/M3/_7_  (.A(a[23]),
    .B(b[23]),
    .Z(\M2/M1/M3/_3_ ));
 OAI21_X1 \M2/M1/M3/_8_  (.A(\M2/M1/M3/_1_ ),
    .B1(\M2/M1/M3/_2_ ),
    .B2(\M2/M1/M3/_0_ ),
    .ZN(c3));
 XNOR2_X1 \M2/M1/M3/_9_  (.A(\M2/M1/M3/_0_ ),
    .B(\M2/M1/M3/_3_ ),
    .ZN(sum[23]));
 INV_X1 \M3/M0/M0/_4_  (.A(c3),
    .ZN(\M3/M0/M0/_0_ ));
 NAND2_X1 \M3/M0/M0/_5_  (.A1(a[24]),
    .A2(b[24]),
    .ZN(\M3/M0/M0/_1_ ));
 NOR2_X1 \M3/M0/M0/_6_  (.A1(a[24]),
    .A2(b[24]),
    .ZN(\M3/M0/M0/_2_ ));
 XOR2_X1 \M3/M0/M0/_7_  (.A(a[24]),
    .B(b[24]),
    .Z(\M3/M0/M0/_3_ ));
 OAI21_X1 \M3/M0/M0/_8_  (.A(\M3/M0/M0/_1_ ),
    .B1(\M3/M0/M0/_2_ ),
    .B2(\M3/M0/M0/_0_ ),
    .ZN(\M3/M0/c1 ));
 XNOR2_X1 \M3/M0/M0/_9_  (.A(\M3/M0/M0/_0_ ),
    .B(\M3/M0/M0/_3_ ),
    .ZN(sum[24]));
 INV_X1 \M3/M0/M1/_4_  (.A(\M3/M0/c1 ),
    .ZN(\M3/M0/M1/_0_ ));
 NAND2_X1 \M3/M0/M1/_5_  (.A1(a[25]),
    .A2(b[25]),
    .ZN(\M3/M0/M1/_1_ ));
 NOR2_X1 \M3/M0/M1/_6_  (.A1(a[25]),
    .A2(b[25]),
    .ZN(\M3/M0/M1/_2_ ));
 XOR2_X1 \M3/M0/M1/_7_  (.A(a[25]),
    .B(b[25]),
    .Z(\M3/M0/M1/_3_ ));
 OAI21_X1 \M3/M0/M1/_8_  (.A(\M3/M0/M1/_1_ ),
    .B1(\M3/M0/M1/_2_ ),
    .B2(\M3/M0/M1/_0_ ),
    .ZN(\M3/M0/c2 ));
 XNOR2_X1 \M3/M0/M1/_9_  (.A(\M3/M0/M1/_0_ ),
    .B(\M3/M0/M1/_3_ ),
    .ZN(sum[25]));
 INV_X1 \M3/M0/M2/_4_  (.A(\M3/M0/c2 ),
    .ZN(\M3/M0/M2/_0_ ));
 NAND2_X1 \M3/M0/M2/_5_  (.A1(a[26]),
    .A2(b[26]),
    .ZN(\M3/M0/M2/_1_ ));
 NOR2_X1 \M3/M0/M2/_6_  (.A1(a[26]),
    .A2(b[26]),
    .ZN(\M3/M0/M2/_2_ ));
 XOR2_X1 \M3/M0/M2/_7_  (.A(a[26]),
    .B(b[26]),
    .Z(\M3/M0/M2/_3_ ));
 OAI21_X1 \M3/M0/M2/_8_  (.A(\M3/M0/M2/_1_ ),
    .B1(\M3/M0/M2/_2_ ),
    .B2(\M3/M0/M2/_0_ ),
    .ZN(\M3/M0/c3 ));
 XNOR2_X1 \M3/M0/M2/_9_  (.A(\M3/M0/M2/_0_ ),
    .B(\M3/M0/M2/_3_ ),
    .ZN(sum[26]));
 INV_X1 \M3/M0/M3/_4_  (.A(\M3/M0/c3 ),
    .ZN(\M3/M0/M3/_0_ ));
 NAND2_X1 \M3/M0/M3/_5_  (.A1(a[27]),
    .A2(b[27]),
    .ZN(\M3/M0/M3/_1_ ));
 NOR2_X1 \M3/M0/M3/_6_  (.A1(a[27]),
    .A2(b[27]),
    .ZN(\M3/M0/M3/_2_ ));
 XOR2_X1 \M3/M0/M3/_7_  (.A(a[27]),
    .B(b[27]),
    .Z(\M3/M0/M3/_3_ ));
 OAI21_X1 \M3/M0/M3/_8_  (.A(\M3/M0/M3/_1_ ),
    .B1(\M3/M0/M3/_2_ ),
    .B2(\M3/M0/M3/_0_ ),
    .ZN(\M3/c1 ));
 XNOR2_X1 \M3/M0/M3/_9_  (.A(\M3/M0/M3/_0_ ),
    .B(\M3/M0/M3/_3_ ),
    .ZN(sum[27]));
 INV_X1 \M3/M1/M0/_4_  (.A(\M3/c1 ),
    .ZN(\M3/M1/M0/_0_ ));
 NAND2_X1 \M3/M1/M0/_5_  (.A1(a[28]),
    .A2(b[28]),
    .ZN(\M3/M1/M0/_1_ ));
 NOR2_X1 \M3/M1/M0/_6_  (.A1(a[28]),
    .A2(b[28]),
    .ZN(\M3/M1/M0/_2_ ));
 XOR2_X1 \M3/M1/M0/_7_  (.A(a[28]),
    .B(b[28]),
    .Z(\M3/M1/M0/_3_ ));
 OAI21_X1 \M3/M1/M0/_8_  (.A(\M3/M1/M0/_1_ ),
    .B1(\M3/M1/M0/_2_ ),
    .B2(\M3/M1/M0/_0_ ),
    .ZN(\M3/M1/c1 ));
 XNOR2_X1 \M3/M1/M0/_9_  (.A(\M3/M1/M0/_0_ ),
    .B(\M3/M1/M0/_3_ ),
    .ZN(sum[28]));
 INV_X1 \M3/M1/M1/_4_  (.A(\M3/M1/c1 ),
    .ZN(\M3/M1/M1/_0_ ));
 NAND2_X1 \M3/M1/M1/_5_  (.A1(a[29]),
    .A2(b[29]),
    .ZN(\M3/M1/M1/_1_ ));
 NOR2_X1 \M3/M1/M1/_6_  (.A1(a[29]),
    .A2(b[29]),
    .ZN(\M3/M1/M1/_2_ ));
 XOR2_X1 \M3/M1/M1/_7_  (.A(a[29]),
    .B(b[29]),
    .Z(\M3/M1/M1/_3_ ));
 OAI21_X1 \M3/M1/M1/_8_  (.A(\M3/M1/M1/_1_ ),
    .B1(\M3/M1/M1/_2_ ),
    .B2(\M3/M1/M1/_0_ ),
    .ZN(\M3/M1/c2 ));
 XNOR2_X1 \M3/M1/M1/_9_  (.A(\M3/M1/M1/_0_ ),
    .B(\M3/M1/M1/_3_ ),
    .ZN(sum[29]));
 INV_X1 \M3/M1/M2/_4_  (.A(\M3/M1/c2 ),
    .ZN(\M3/M1/M2/_0_ ));
 NAND2_X1 \M3/M1/M2/_5_  (.A1(a[30]),
    .A2(b[30]),
    .ZN(\M3/M1/M2/_1_ ));
 NOR2_X1 \M3/M1/M2/_6_  (.A1(a[30]),
    .A2(b[30]),
    .ZN(\M3/M1/M2/_2_ ));
 XOR2_X1 \M3/M1/M2/_7_  (.A(a[30]),
    .B(b[30]),
    .Z(\M3/M1/M2/_3_ ));
 OAI21_X1 \M3/M1/M2/_8_  (.A(\M3/M1/M2/_1_ ),
    .B1(\M3/M1/M2/_2_ ),
    .B2(\M3/M1/M2/_0_ ),
    .ZN(\M3/M1/c3 ));
 XNOR2_X1 \M3/M1/M2/_9_  (.A(\M3/M1/M2/_0_ ),
    .B(\M3/M1/M2/_3_ ),
    .ZN(sum[30]));
 INV_X1 \M3/M1/M3/_4_  (.A(\M3/M1/c3 ),
    .ZN(\M3/M1/M3/_0_ ));
 NAND2_X1 \M3/M1/M3/_5_  (.A1(a[31]),
    .A2(b[31]),
    .ZN(\M3/M1/M3/_1_ ));
 NOR2_X1 \M3/M1/M3/_6_  (.A1(a[31]),
    .A2(b[31]),
    .ZN(\M3/M1/M3/_2_ ));
 XOR2_X1 \M3/M1/M3/_7_  (.A(a[31]),
    .B(b[31]),
    .Z(\M3/M1/M3/_3_ ));
 OAI21_X1 \M3/M1/M3/_8_  (.A(\M3/M1/M3/_1_ ),
    .B1(\M3/M1/M3/_2_ ),
    .B2(\M3/M1/M3/_0_ ),
    .ZN(cout));
 XNOR2_X1 \M3/M1/M3/_9_  (.A(\M3/M1/M3/_0_ ),
    .B(\M3/M1/M3/_3_ ),
    .ZN(sum[31]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_113 ();
endmodule
